---------------------------------------------------------------------------------
-- This is free and unencumbered software released into the public domain.
--
-- Anyone is free to copy, modify, publish, use, compile, sell, or
-- distribute this software, either in source code form or as a compiled
-- binary, for any purpose, commercial or non-commercial, and by any
-- means.
--
-- In jurisdictions that recognize copyright laws, the author or authors
-- of this software dedicate any and all copyright interest in the
-- software to the public domain. We make this dedication for the benefit
-- of the public at large and to the detriment of our heirs and
-- successors. We intend this dedication to be an overt act of
-- relinquishment in perpetuity of all present and future rights to this
-- software under copyright law.
--
-- THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
-- EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
-- MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT.
-- IN NO EVENT SHALL THE AUTHORS BE LIABLE FOR ANY CLAIM, DAMAGES OR
-- OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE,
-- ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR
-- OTHER DEALINGS IN THE SOFTWARE.
--
-- For more information, please refer to <http://unlicense.org/>
---------------------------------------------------------------------------------


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity rom_128x10_exclif2_ip is
    port (
        clka : in std_logic;
        addra : in std_logic_vector(6 downto 0);
        douta : out std_logic_vector(39 downto 0)
    );
end entity rom_128x10_exclif2_ip;

architecture behavior of rom_128x10_exclif2_ip is


    type rom_type is array (0 to 128) of std_logic_vector(39 downto 0);


    constant mem : rom_type := (
"0000000000000000000000001111000000001111",
"0000111100000000000011110000000000000001",
"0000000000000000000000000000000011110000",
"0000000000000001000000000000000000000000",
"0000000000000000000000011111000000000000",
"0000000011111111111100000000000011110000",
"0000000000000000000000000000000000001111",
"0000000100000000000100000000000000000000",
"0001000000010001000000000000000100000000",
"0000000011110000000100000000111100001111",
"0000000000000000000000001111000000000001",
"0001000100010000000100000000000000010000",
"1111000011110000000000000001000000000001",
"0000111100000000000000010000000000000000",
"0000000100000000000000000000000100010000",
"0000000011110001000000000000000100000000",
"0000000000000000000000001111000100000000",
"0000111100000000000000001111000000001111",
"0000000011110000111100000000000000010000",
"1111000000000000000000000000111111110000",
"0000000000000000000000000000000000000000",
"1111000011110000000011110000000000000000",
"0000000000000000111100001111000011110000",
"0000000000000000000000000000000000010000",
"1111000000000000000000000000000000000000",
"0000000000000000000000001111000000000000",
"0000000000000000000000010000111100000000",
"0001000100010000000000000000000011111111",
"0000000011110000000011110000000100010000",
"0000000000001111000000000000000000000000",
"0000000000000000000000010000000111111111",
"0001000000000000000100000000000000000000",
"0000111100000000111100000001000000000000",
"0000000000000000000000001111000100000001",
"0000000000000000000000000000000011111111",
"0000000000000000000100000001000011110001",
"0000000111111111000000000000000000000000",
"0000000100000000000000000000000000000000",
"0000000100000000000000000000000011110000",
"0000111100010000000000000000000000001111",
"0000000000000001000000000000000000000000",
"0000000000010000000000000001000000000000",
"1111000000000000000000011111111100000000",
"0000000000010000000000011111000011110000",
"0000000000000001111100000000000011110000",
"0000000011110000000000000001000000000000",
"0000000000000001111100001111000000000000",
"0000111100000000000011110001111100000000",
"0000000000001111000000000000111111110000",
"1111000000010000000000000000000000001111",
"1111000100000000000000000000000000000000",
"1111000000000001000100000001000000000000",
"0000000000000001111100000000000000000000",
"0000000000000001111111110000000000000000",
"0000000000001111111111110000000011111111",
"0000000000000000000000000000000011110000",
"0000000000001111000100000000000000000000",
"0000000000000000111100000000111111111111",
"1111000000000000000000000000111100000000",
"0000000100000000000000000000111111111111",
"0000000000000001000000000001000000010000",
"0000000011110000000000000000000100000000",
"0000000000010001000000000000000000001111",
"0000000000000000111100000000000000000000",
"0001000011110000000000000000000000000000",
"1111000100000000000100000000111100000000",
"1111111100000000111100010000000011110001",
"0000000000000001000100000000000000000000",
"0000000100000000111100000000000000000000",
"0001000011110000000000000000000000000000",
"0000000000000000000000000000000000001111",
"1111000011110000111100000001000011110000",
"0000111100000000000011110000000111110001",
"0000000100000000000011110000000000000001",
"0000000000000000000000000000000011110000",
"0000000000001111000011111111111100000000",
"0000000100000000000000000000111100010000",
"0000000100000000111100000001000011110000",
"0001000100000000111100001111000100000000",
"0001000000000000000000001111000000000000",
"0000000000000000000100000000000000000000",
"0000111100000000111100001111000000010001",
"1111000000000001000000000000000000000000",
"1111000011110000000000000000000000000000",
"1111000000010000111111110001111100000001",
"0000000000000000000000000000000100000001",
"0000000100001111000100000000000100000001",
"0000000000000000000000010000000000000000",
"1111000000010001000100010000000000000000",
"0000000000010001000000001111000000000000",
"0000000011110001111111110000000011110000",
"1111000000001111000000001111000100000000",
"0000000000000000000000000000000000000000",
"0000000000000001000000000000000000000000",
"0000000100000000111100000000000000000000",
"0000000000010000111100001111111100000000",
"0001000000000001000000000000111100000000",
"0000111100000000000000001111000000010000",
"0000111100000000000000000000000011110000",
"0000000000011111000000010001000000000000",
"0001000000001111111100000001000000010000",
"0000000000000000000000000000000000000000",
"0000000011110000000011110000000000000001",
"0000000011110000000000010000000000000000",
"1111000000001111000000001111000000010000",
"0000000000000000000000010000000000000000",
"1111000011110000000000000001000011110001",
"1111000100000000000000001111000100000000",
"0000000000000000000100000000000100000000",
"1111111100000000000011110000000000000000",
"0000111111111111000000001111000111110000",
"0000000000001111000000010000000000000000",
"0000000000010000000000000000000000010001",
"0001000000001111000000010000000000000001",
"0000000000000000000011110000111100000000",
"0000000000000000000000000000000000001111",
"0001111111110000000000000000000000000000",
"0000000000000000000000001111000100000000",
"0000000100000001000000000000000000001111",
"0000000000010000000000001111000000010000",
"0000000000000001111100000000111111110001",
"0001000000000000111100000001111100000000",
"0001000000000000000000001111000100010000",
"0000000000001111000000001111000000001111",
"0001000100010001000000000001000100000000",
"0000000100001111000000000000000011110000",
"0000000100011111000000000000000000000000",
"0000000011110000000000000001111111110001",
"0000000000000000000000000000000000000000");

begin

    rom_behavior : process(clka )
    begin

        if clka'event and clka='1' 
        then

            douta <= mem(to_integer(unsigned(addra)));

        end if;

    end process rom_behavior;


end architecture behavior;

